library verilog;
use verilog.vl_types.all;
entity akkumulator_vlg_vec_tst is
end akkumulator_vlg_vec_tst;
